19/09/2019 10:29:08:GuestPageNew.aspx :: Page_Load ::    at System.Data.DataRow.GetDataColumn(String columnName)
   at System.Data.DataRow.get_Item(String columnName)
   at GuestPagenew.BindFlightDetailsAmend() in D:\AgentsOnline_New\GuestPagenew.aspx.vb:line 1422
   at GuestPagenew.LoadHome() in D:\AgentsOnline_New\GuestPagenew.aspx.vb:line 606
   at GuestPagenew.Page_Load(Object sender, EventArgs e) in D:\AgentsOnline_New\GuestPagenew.aspx.vb:line 68:: admin
19/09/2019 10:29:23:GuestPageNew.aspx :: Page_Load ::    at System.Data.DataRow.GetDataColumn(String columnName)
   at System.Data.DataRow.get_Item(String columnName)
   at GuestPagenew.BindFlightDetailsAmend() in D:\AgentsOnline_New\GuestPagenew.aspx.vb:line 1422
   at GuestPagenew.LoadHome() in D:\AgentsOnline_New\GuestPagenew.aspx.vb:line 606
   at GuestPagenew.Page_Load(Object sender, EventArgs e) in D:\AgentsOnline_New\GuestPagenew.aspx.vb:line 68:: admin
19/09/2019 10:34:29:GuestPageNew.aspx :: Page_Load ::    at System.Data.DataRow.GetDataColumn(String columnName)
   at System.Data.DataRow.get_Item(String columnName)
   at GuestPagenew.BindFlightDetailsAmend() in D:\AgentsOnline_New\GuestPagenew.aspx.vb:line 1422
   at GuestPagenew.LoadHome() in D:\AgentsOnline_New\GuestPagenew.aspx.vb:line 606
   at GuestPagenew.Page_Load(Object sender, EventArgs e) in D:\AgentsOnline_New\GuestPagenew.aspx.vb:line 68:: admin
19/09/2019 10:36:52:GuestPageNew.aspx :: Page_Load ::    at System.Data.DataRow.GetDataColumn(String columnName)
   at System.Data.DataRow.get_Item(String columnName)
   at GuestPagenew.BindFlightDetailsAmend() in D:\AgentsOnline_New\GuestPagenew.aspx.vb:line 1453
   at GuestPagenew.LoadHome() in D:\AgentsOnline_New\GuestPagenew.aspx.vb:line 606
   at GuestPagenew.Page_Load(Object sender, EventArgs e) in D:\AgentsOnline_New\GuestPagenew.aspx.vb:line 68:: admin
19/09/2019 13:02:39:Login.aspx:: GetIpLocationName :: The remote server returned an error: (403) Forbidden.
19/09/2019 13:02:56:MyAccount.aspx :: lbEdit_Click :: Thread was being aborted.:: admin
19/09/2019 13:13:57:GuestPageNew.aspx :: Page_Load ::    at System.Threading.Thread.AbortInternal()
   at System.Threading.Thread.Abort(Object stateInfo)
   at System.Web.HttpResponse.AbortCurrentThread()
   at System.Web.HttpResponse.End()
   at System.Web.HttpResponse.Redirect(String url, Boolean endResponse, Boolean permanent)
   at System.Web.HttpResponse.Redirect(String url, Boolean endResponse)
   at GuestPagenew.Page_Load(Object sender, EventArgs e) in D:\AgentsOnline_New\GuestPagenew.aspx.vb:line 36:: 
19/09/2019 13:14:04:Login.aspx:: GetIpLocationName :: The remote server returned an error: (403) Forbidden.
19/09/2019 13:14:26:MyAccount.aspx :: lbEdit_Click :: Thread was being aborted.:: admin
19/09/2019 13:40:11:MyAccount.aspx :: lbEdit_Click :: Thread was being aborted.:: admin
19/09/2019 13:50:27:MyAccount.aspx :: lbEdit_Click :: Thread was being aborted.:: admin
19/09/2019 15:10:42:Login.aspx:: GetIpLocationName :: The remote server returned an error: (403) Forbidden.
19/09/2019 15:11:45:HotelSearch.aspx :: btnBookNow_Click :: Thread was being aborted.:: admin
19/09/2019 15:12:25:HotelSearch.aspx :: btnBookNow_Click :: Thread was being aborted.:: admin
19/09/2019 15:13:21:AirportMeetSearch.aspx :: btnBookNow_Click :: Thread was being aborted.:: admin
19/09/2019 15:13:43:TransferSearch.aspx :: btnBookNow_Click :: Thread was being aborted.:: admin
19/09/2019 15:16:03:HotelSearch.aspx :: btnBookNow_Click :: Thread was being aborted.:: admin
19/09/2019 16:38:25:MyAccount.aspx :: lbEdit_Click :: Thread was being aborted.:: admin
19/09/2019 16:59:00:Login.aspx:: GetIpLocationName :: The remote server returned an error: (403) Forbidden.
19/09/2019 16:59:24:Invalid object name 'priceadults'. :: GetDataSet
19/09/2019 16:59:44:Invalid object name 'priceadults'. :: GetDataSet
19/09/2019 17:00:31:Invalid object name 'priceadults'. :: GetDataSet
19/09/2019 17:00:32:HotelSearch.aspx :: btnPreHotelSave_Click :: Object reference not set to an instance of an object.:: admin
19/09/2019 17:00:58:Login.aspx:: GetIpLocationName :: The remote server returned an error: (403) Forbidden.
19/09/2019 17:02:09:HotelSearch.aspx :: btnBookNow_Click :: Thread was being aborted.:: admin
19/09/2019 17:02:28:Invalid object name 'priceadults'. :: GetDataSet
19/09/2019 17:02:50:Invalid object name 'priceadults'. :: GetDataSet
19/09/2019 17:03:00:Invalid object name 'priceadults'. :: GetDataSet
19/09/2019 17:03:16:Invalid object name 'priceadults'. :: GetDataSet
19/09/2019 17:03:49:HotelSearch.aspx :: btnBookNow_Click :: Thread was being aborted.:: admin
19/09/2019 17:09:19:HotelSearch.aspx :: btnBookNow_Click :: Thread was being aborted.:: admin
19/09/2019 17:44:11:Login.aspx:: GetIpLocationName :: The remote server returned an error: (403) Forbidden.
19/09/2019 17:44:28:Invalid object name 'priceadults'. :: GetDataSet
19/09/2019 17:44:49:HotelSearch.aspx :: btnBookNow_Click :: Thread was being aborted.:: admin
19/09/2019 17:45:27:HotelSearch.aspx :: btnBookNow_Click :: Thread was being aborted.:: admin
19/09/2019 17:46:08:HotelSearch.aspx :: btnBookNow_Click :: Thread was being aborted.:: admin
19/09/2019 17:48:24:HotelSearch.aspx :: btnBookNow_Click :: Thread was being aborted.:: admin
19/09/2019 18:58:22:MyAccount.aspx :: lbEdit_Click :: Thread was being aborted.:: admin
19/09/2019 19:13:38:Login.aspx:: GetIpLocationName :: The remote server returned an error: (403) Forbidden.
19/09/2019 19:15:29:   at System.Data.SqlClient.SqlConnection.OnError(SqlException exception, Boolean breakConnection, Action`1 wrapCloseInAction)
   at System.Data.SqlClient.SqlInternalConnection.OnError(SqlException exception, Boolean breakConnection, Action`1 wrapCloseInAction)
   at System.Data.SqlClient.TdsParser.ThrowExceptionAndWarning(TdsParserStateObject stateObj, Boolean callerHasConnectionLock, Boolean asyncClose)
   at System.Data.SqlClient.TdsParser.TryRun(RunBehavior runBehavior, SqlCommand cmdHandler, SqlDataReader dataStream, BulkCopySimpleResultSet bulkCopyHandler, TdsParserStateObject stateObj, Boolean& dataReady)
   at System.Data.SqlClient.SqlCommand.FinishExecuteReader(SqlDataReader ds, RunBehavior runBehavior, String resetOptionsString, Boolean isInternal, Boolean forDescribeParameterEncryption, Boolean shouldCacheForAlwaysEncrypted)
   at System.Data.SqlClient.SqlCommand.RunExecuteReaderTds(CommandBehavior cmdBehavior, RunBehavior runBehavior, Boolean returnStream, Boolean async, Int32 timeout, Task& task, Boolean asyncWrite, Boolean inRetry, SqlDataReader ds, Boolean describeParameterEncryptionRequest)
   at System.Data.SqlClient.SqlCommand.RunExecuteReader(CommandBehavior cmdBehavior, RunBehavior runBehavior, Boolean returnStream, String method, TaskCompletionSource`1 completion, Int32 timeout, Task& task, Boolean& usedCache, Boolean asyncWrite, Boolean inRetry)
   at System.Data.SqlClient.SqlCommand.InternalExecuteNonQuery(TaskCompletionSource`1 completion, String methodName, Boolean sendToPipe, Int32 timeout, Boolean& usedCache, Boolean asyncWrite, Boolean inRetry)
   at System.Data.SqlClient.SqlCommand.ExecuteNonQuery()
   at clsUtilities.ExecuteNonQuery_Param(String storedProcedure, List`1 sqlParamList) in D:\AgentsOnline_New\App_Code\DAL\clsUtilities.vb:line 549 :: ExecuteNonQuery_Param
19/09/2019 19:15:29:MyAccount.aspx :: lbQEdit_Click :: Thread was being aborted.:: admin
19/09/2019 19:16:10:   at System.Data.SqlClient.SqlConnection.OnError(SqlException exception, Boolean breakConnection, Action`1 wrapCloseInAction)
   at System.Data.SqlClient.SqlInternalConnection.OnError(SqlException exception, Boolean breakConnection, Action`1 wrapCloseInAction)
   at System.Data.SqlClient.TdsParser.ThrowExceptionAndWarning(TdsParserStateObject stateObj, Boolean callerHasConnectionLock, Boolean asyncClose)
   at System.Data.SqlClient.TdsParser.TryRun(RunBehavior runBehavior, SqlCommand cmdHandler, SqlDataReader dataStream, BulkCopySimpleResultSet bulkCopyHandler, TdsParserStateObject stateObj, Boolean& dataReady)
   at System.Data.SqlClient.SqlCommand.FinishExecuteReader(SqlDataReader ds, RunBehavior runBehavior, String resetOptionsString, Boolean isInternal, Boolean forDescribeParameterEncryption, Boolean shouldCacheForAlwaysEncrypted)
   at System.Data.SqlClient.SqlCommand.RunExecuteReaderTds(CommandBehavior cmdBehavior, RunBehavior runBehavior, Boolean returnStream, Boolean async, Int32 timeout, Task& task, Boolean asyncWrite, Boolean inRetry, SqlDataReader ds, Boolean describeParameterEncryptionRequest)
   at System.Data.SqlClient.SqlCommand.RunExecuteReader(CommandBehavior cmdBehavior, RunBehavior runBehavior, Boolean returnStream, String method, TaskCompletionSource`1 completion, Int32 timeout, Task& task, Boolean& usedCache, Boolean asyncWrite, Boolean inRetry)
   at System.Data.SqlClient.SqlCommand.InternalExecuteNonQuery(TaskCompletionSource`1 completion, String methodName, Boolean sendToPipe, Int32 timeout, Boolean& usedCache, Boolean asyncWrite, Boolean inRetry)
   at System.Data.SqlClient.SqlCommand.ExecuteNonQuery()
   at clsUtilities.ExecuteNonQuery_Param(String storedProcedure, List`1 sqlParamList) in D:\AgentsOnline_New\App_Code\DAL\clsUtilities.vb:line 549 :: ExecuteNonQuery_Param
19/09/2019 19:16:10:MyAccount.aspx :: lbQEdit_Click :: Thread was being aborted.:: admin
